module rom_instructions
#(parameter DATA_WIDTH=32, parameter ADDR_WIDTH=32, parameter ROM_SIZE = 800)
(
	input [(ADDR_WIDTH-1):0] addr,
	input clk, 
	output reg [(DATA_WIDTH-1):0] q
);

	 // Ajuste do tamanho do vetor ROM
    reg [DATA_WIDTH-1:0] rom [0:ROM_SIZE-1];

    // Indexação limitada para evitar endereços inválidos
    wire [$clog2(ROM_SIZE)-1:0] addr_index = addr[$clog2(ROM_SIZE)-1:0];

	// Initialize the ROM with $readmemb.  Put the memory contents
	// in the file single_port_rom_init.txt.  Without this file,
	// this design will not compile.

	// See Verilog LRM 1364-2001 Section 17.2.8 for details on the
	// format of this file, or see the "Using $readmemb and $readmemh"
	// template later in this section.

	initial
	begin
		//rotina
			$readmemb("instrucoes_ram/rotina_troca_contexto.txt", rom, 0, 199);
			//sistema operacional
			$readmemb("instrucoes_ram/so.txt", rom, 200, 399);
			//soma
			$readmemb("instrucoes_ram/programa_1.txt", rom, 400, 599);
			//subtracao
			$readmemb("instrucoes_ram/programa_2.txt", rom, 600, 799);
			//maior
			//$readmemb("instrucoes_ram/programa_3.txt", rom, 800, 999);
			//fibonacci
			//$readmemb("instrucoes_ram/programa_4.txt", rom, 1000, 1199);
			//perimetro
			//$readmemb("instrucoes_ram/programa_5.txt", rom, 1200, 1399);
			//gcd
			//$readmemb("instrucoes_ram/programa_6.txt", rom, 1400, 1599);
			//fatorial
			//$readmemb("instrucoes_ram/programa_7.txt", rom, 1600, 1799);
			//potencia
			//$readmemb("instrucoes_ram/programa_8.txt", rom, 1800, 1999);
	end

	always_ff @(posedge clk)
	begin
		q <= rom[addr];
	end

endmodule
