module game_process (
input clock,
output );
endmodule 