module display7seg (input[31:0] segmentos, input[31:0] segmentosPrograma, input neg, output reg[6:0] seg[7:0]);

	
	always @ (*) begin
		case (segmentos[3:0])
			4'b0000: seg[0] = 7'b1000000;
			4'b0001: seg[0] = 7'b1111001;
			4'b0010: seg[0] = 7'b0100100;
			4'b0011: seg[0] = 7'b0110000;
			4'b0100: seg[0] = 7'b0011001;
			4'b0101: seg[0] = 7'b0010010;
			4'b0110: seg[0] = 7'b0000010;
			4'b0111: seg[0] = 7'b1111000;
			4'b1000: seg[0] = 7'b0000000;
			4'b1001: seg[0] = 7'b0011000;
			default: seg[0] = 7'b1111111;
		endcase
		case (segmentos[7:4])
			4'b0000: seg[1] = 7'b1000000;
			4'b0001: seg[1] = 7'b1111001;
			4'b0010: seg[1] = 7'b0100100;
			4'b0011: seg[1] = 7'b0110000;
			4'b0100: seg[1] = 7'b0011001;
			4'b0101: seg[1] = 7'b0010010;
			4'b0110: seg[1] = 7'b0000010;
			4'b0111: seg[1] = 7'b1111000;
			4'b1000: seg[1] = 7'b0000000;
			4'b1001: seg[1] = 7'b0011000;
			default: seg[1] = 7'b1111111;
		endcase
		case (segmentos[11:8])
			4'b0000: seg[2] = 7'b1000000;
			4'b0001: seg[2] = 7'b1111001;
			4'b0010: seg[2] = 7'b0100100;
			4'b0011: seg[2] = 7'b0110000;
			4'b0100: seg[2] = 7'b0011001;
			4'b0101: seg[2] = 7'b0010010;
			4'b0110: seg[2] = 7'b0000010;
			4'b0111: seg[2] = 7'b1111000;
			4'b1000: seg[2] = 7'b0000000;
			4'b1001: seg[2] = 7'b0011000;
			default: seg[2] = 7'b1111111;
		endcase
		case (segmentos[15:12])
			4'b0000: seg[3] = 7'b1000000;
			4'b0001: seg[3] = 7'b1111001;
			4'b0010: seg[3] = 7'b0100100;
			4'b0011: seg[3] = 7'b0110000;
			4'b0100: seg[3] = 7'b0011001;
			4'b0101: seg[3] = 7'b0010010;
			4'b0110: seg[3] = 7'b0000010;
			4'b0111: seg[3] = 7'b1111000;
			4'b1000: seg[3] = 7'b0000000;
			4'b1001: seg[3] = 7'b0011000;
			default: seg[3] = 7'b1111111;
		endcase
		case (segmentos[19:16])
			4'b0000: seg[4] = 7'b1000000;
			4'b0001: seg[4] = 7'b1111001;
			4'b0010: seg[4] = 7'b0100100;
			4'b0011: seg[4] = 7'b0110000;
			4'b0100: seg[4] = 7'b0011001;
			4'b0101: seg[4] = 7'b0010010;
			4'b0110: seg[4] = 7'b0000010;
			4'b0111: seg[4] = 7'b1111000;
			4'b1000: seg[4] = 7'b0000000;
			4'b1001: seg[4] = 7'b0011000;
			default: seg[4] = 7'b1111111;
		endcase
		case (segmentos[23:20])
			4'b0000: seg[5] = 7'b1000000;
			4'b0001: seg[5] = 7'b1111001;
			4'b0010: seg[5] = 7'b0100100;
			4'b0011: seg[5] = 7'b0110000;
			4'b0100: seg[5] = 7'b0011001;
			4'b0101: seg[5] = 7'b0010010;
			4'b0110: seg[5] = 7'b0000010;
			4'b0111: seg[5] = 7'b1111000;
			4'b1000: seg[5] = 7'b0000000;
			4'b1001: seg[5] = 7'b0011000;
			default: seg[5] = 7'b1111111;
		endcase
		case ({segmentosPrograma[15:12], segmentosPrograma[11:8]})
			 8'b00000000, 8'b00000001: begin
				  seg[7] = 7'b1111111; 
				  seg[6] = 7'b1000000; // 0
			 end
			 8'b00000010, 8'b00000011: begin
				  seg[7] = 7'b1111111;
				  seg[6] = 7'b1000000; // 0
			 end
			 8'b00000100, 8'b00000101: begin
				  seg[7] = 7'b1111111;
				  seg[6] = 7'b1111001; // 1
			 end
			 8'b00000110, 8'b00000111: begin
				  seg[7] = 7'b1111111;
				  seg[6] = 7'b0100100; // 2
			 end
			 8'b00001000, 8'b00001001: begin
				  seg[7] = 7'b1111111;
				  seg[6] = 7'b0110000; // 3
			 end
			 8'b00010000, 8'b00010001: begin
				  seg[7] = 7'b1111111;
				  seg[6] = 7'b0011001; // 4
			 end
			 8'b00010010, 8'b00010011: begin
				  seg[7] = 7'b1111111;
				  seg[6] = 7'b0010010; // 5
			 end
			 8'b00010100, 8'b00010101: begin
				  seg[7] = 7'b1111111;
				  seg[6] = 7'b0000010; // 6
			 end
			 8'b00010110, 8'b00010111: begin
				  seg[7] = 7'b1111111;
				  seg[6] = 7'b1111000; // 7
			 end
			 8'b00011000, 8'b00011001: begin
				  seg[7] = 7'b1111111;
				  seg[6] = 7'b0000000; // 8
			 end
			 default: begin
				  seg[7] = 7'b1111111;
				  seg[6] = 7'b1111111; // Caso inválido
			 end
		endcase
		if(neg)begin
		seg[7] = 7'b0111111;
		end
	end
endmodule
		